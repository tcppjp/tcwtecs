/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

/**
 * TCWTecs infrastructure. Do not call any members in the user application.
 */
signature sTWTimerLink {
};
