/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("sTWDispatchTarget.cdl");
import("TWTypes.cdl");

signature sTWDispatcherControl {
    /**
     * ディスパッチターゲットと引数を指定して、呼出しを行います。
     *
     * ターゲットは、指定された引数を使用して、GUIスレッドで呼び出されます。
     * 本関数の呼出しは、ターゲットの呼出しが完了した後に返ります。
     *
     * 本関数によるディスパッチは同期的であり、従って割込みハンドラ等では使用できません。
     * 割込みハンドラからディスパッチを行う場合、tTWDeferredDispatch を使用してください。
     */
    void invoke([in] Descriptor(sTWDispatchTarget) target, [in] intptr_t param);

    /**
     * 時刻を取得します。基準とする時刻は任意ですが、それは変化しません。取得される時刻は stable です。
     */
    TWTimePoint getTime(void);
};
