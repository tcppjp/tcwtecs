/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTecs.cdl");
import("tTWSDLDispatcher.cdl");
import("tTWSDLGraphicsDevice.cdl");

import("tSimpleButton.cdl");
import("tSDLApp.cdl");

cell tTWSDLDispatcher Dispatcher {
};

cell tTWTimerManager TimerManager {
	cDispatcherLink = Dispatcher.eDispatcherLink;
	eTimerManager <= Dispatcher.cTimerManager;
};

cell tTWKeyboardInputManager KeyboardInputManager {
};

cell tTWTouchInputManager TouchInputManager {
	maxNumTouches = 1;
	cElement[0] = TouchInputManager.eNullElementLink;
};

cell tTWSDLGraphicsDevice SDL {
	width = 120;
	height = 120;
	title = "Hello World!";
	windowFlags = C_EXP("0");

	eSDLEvent <= Dispatcher.cSDLEvent[0];

	cKeyboardInputDriverEvent = KeyboardInputManager.eDriverEvent;
	cTouchInputDriverEvent = TouchInputManager.eDriverEvent;
};

cell tTWDesktop Desktop {
	cGraphicsDevice = SDL.eGraphicsDevice;
	eGraphicsDevice <= SDL.cGraphicsDevice;
	cTimerManager = TimerManager.eTimerManager;
};

celltype tMainWindowCore {
	entry sTWPaintEvent ePaintEvent;
	call sTWDrawingContext cDC;

	entry sAction eButtonActivated[3];
};

composite tMainWindow {
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;
	call sTWDesktopLink cDesktopLink;

	entry sTWTouchInputSubviewLink eTouchInputSuperview;
	call sTWTouchInputSuperviewLink cTouchInputSuperview;

	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	cell tSimpleButton Button1;
	cell tSimpleButton Button2;
	cell tSimpleButton Button3;

	cell tMainWindowCore Core;

	cell tTWStaticRectSource View_Bounds {
		x = 0; y = 0; w = 120; h = 120;
	};
	cell tTWStaticViewStyleSource View_Style {
		value = C_EXP("TWViewStyleVisible");
	};

	cell tTWView View {
		cSuperview => composite.cSuperview;
		cDesktopLink => composite.cDesktopLink;

		cBoundsSource = View_Bounds.eSource;
		cStyleSource = View_Style.eSource;

		// TODO: コールバック結合で記述したい
		cSubview[0] = Button1.eSuperview;
		cSubview[1] = Button2.eSuperview;
		cSubview[2] = Button3.eSuperview;

		cPaintEvent = Core.ePaintEvent;
	};
	composite.eSuperview => View.eSuperview;

	cell tTWTouchInputElement TouchInputElement {
		cSubview[0] = Button1.eTouchInputSuperview;
		cSubview[1] = Button2.eTouchInputSuperview;
		cSubview[2] = Button3.eTouchInputSuperview;

		cSuperview => composite.cTouchInputSuperview;

		cBoundsSource = View_Bounds.eSource;
		cStyleSource = View_Style.eSource;
	};
	composite.eTouchInputSuperview => TouchInputElement.eSuperview;

	cell tMainWindowCore Core {
		cDC = View.eDrawingContext;
	};

	cell tTWStaticRectSource Button1_Bounds {
		x = 20; y = 20; w = 80; h = 20;
	};
	cell tTWStaticRectSource Button2_Bounds {
		x = 20; y = 50; w = 80; h = 20;
	};
	cell tTWStaticRectSource Button3_Bounds {
		x = 20; y = 80; w = 80; h = 20;
	};
	cell tTWStaticViewStyleSource Button_Style {
		value = C_EXP("TWViewStyleVisible");
	};
	cell tSimpleButton Button1 {
		cSuperview = View.eSubview[0];
		cTouchInputSuperview = TouchInputElement.eSubview[0];
		cDesktopLink => composite.cDesktopLink;
		cKeyboardInputManager => composite.cKeyboardInputManager;

		cBoundsSource = Button1_Bounds.eSource;
		cStyleSource = Button_Style.eSource;

		cAction = Core.eButtonActivated[0];
	};
	cell tSimpleButton Button2 {
		cSuperview = View.eSubview[1];
		cTouchInputSuperview = TouchInputElement.eSubview[1];
		cDesktopLink => composite.cDesktopLink;
		cKeyboardInputManager => composite.cKeyboardInputManager;

		cBoundsSource = Button2_Bounds.eSource;
		cStyleSource = Button_Style.eSource;

		cAction = Core.eButtonActivated[1];
	};
	cell tSimpleButton Button3 {
		cSuperview = View.eSubview[2];
		cTouchInputSuperview = TouchInputElement.eSubview[2];
		cDesktopLink => composite.cDesktopLink;
		cKeyboardInputManager => composite.cKeyboardInputManager;

		cBoundsSource = Button3_Bounds.eSource;
		cStyleSource = Button_Style.eSource;

		cAction = Core.eButtonActivated[2];
	};
};

cell tMainWindow MainWindow {
	cSuperview = Desktop.eSubview;
	eSuperview <= Desktop.cSubview;
	cDesktopLink = Desktop.eDesktopLink;
	cKeyboardInputManager = KeyboardInputManager.eControl;

	cTouchInputSuperview = TouchInputManager.eSubview;
	eTouchInputSuperview <= TouchInputManager.cSubview;
};

cell tSDLApp App {
	cSDL = SDL.eControl;
	cSDLDispatcher = Dispatcher.eSDLDispatcher;

	cDesktop = Desktop.eDesktop;
};
