/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");

// import_C("tecsui/colors.h");
// import_C("tecsui/geometry.h");
// import_C("tecsui/bitmap.h");

signature sTWGraphicsDeviceOutput
{
	void getScreenSize([out] TWSize *outSize);
	[oneway] void setClippingRect([in] const TWRect *rect);
	[oneway] void subtractClippingRect([in] const TWRect *rect);
	[oneway] void fillRect([in] TWColor color, [in] const TWRect *rect);
	[oneway] void drawBitmap(
		[in, size_is(numBytes)] const char *data,
		[in] TWPixelFormat format,
		[in] const TWSize *bitmapSize,
		[in] uint32_t numBytes,
		[in] const TWRect *inRect,
		[in] const TWPoint *outLoc,
		[in] TWColor monoColor);
	[oneway] void update([in] const TWRect *rect);
};
