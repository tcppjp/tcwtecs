/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTypes.cdl");

/**
 * TCWTecs infrastructure. Do not call any members in the user application.
 */
[callback]
signature sTWSubviewLink
{
	/**
	 * @param clipRect Region to be updated (in global coordinate)
	 * @param globalBounds Bounding rect of the caller (in global coordinate)
	 */
	void paint([in] const TWRect *clipRect, [in] const TWRect *globalBounds);

    /**
     * @param clipRect Region to be updated (in global coordinate)
     * @param mode 0: no TWViewStyleClipSiblings only, 1: TWViewStyleClipSiblings only
     */
    void subtractClippingRect([in] const TWRect *clipRect, [in] const TWRect *globalBounds, [in] uint8_t mode);
};
