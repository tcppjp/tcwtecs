[callback]
signature sAction {
	void activated(void);
};
