/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");

signature sTWDeferredDispatchControl
{
    /**
     * 遅延ディスパッチをスケジュールします。
     *
     * TODO: should update `param` if it's already active?
     *
     * ディスパッチャがクリティカルセクションに進入した状態でない限り、任意のコンテクストから
     * 呼び出せます。
     *
     * @return 既にスケジュール済みであった場合は 0、それ以外の場合は 1。
     */
    uint8_t start([in] intptr_t param);

    /**
     * 遅延ディスパッチをキャンセルします。
     *
     * ディスパッチャがクリティカルセクションに進入した状態でない限り、任意のコンテクストから
     * 呼び出せます。
     *
     * @return スケジュールされていなかった場合は 0、それ以外の場合は 1。
     */
    uint8_t cancel(void);

    // TODO: join (or wait)?
};
