/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import_C("tecsui/private.h");

/**
 * TCWTecs infrastructure. Do not call any members in the user application.
 */
[deviate, callback]
signature sTWTimerManagerLink {
    /**
     * Called by a timer.
     *
     * Prerequisite: `!(timer->flags & (kTWTimerFlagsActive | kTWTimerFlagsPending))`
     */
    void registerTimer([inout] TWTimerDescriptor *timer);

    /**
     * Called by a timer.
     *
     * Prerequisite: `timer->flags & (kTWTimerFlagsActive | kTWTimerFlagsPending)`
     */
    void unregisterTimer([inout] TWTimerDescriptor *timer);

    /** Called by a deferred dispatch */
    uint8_t registerDeferredDispatch([inout] TWDeferredDispatchDescriptor *dd, [in] intptr_t param);

    /** Called by a deferred dispatch */
    uint8_t unregisterDeferredDispatch([inout] TWDeferredDispatchDescriptor *dd);

    /** Called by a dispatcher */
    void handleTimeout(void);

    /** Called by a dispatcher */
    void handleDeferredDispatch(void);
};
