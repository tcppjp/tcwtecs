/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("sTWDispatcherControl.cdl");
import("sTWDispatchTarget.cdl");
import("sTWDispatcherLink.cdl");
import("sTWTimerManagerLink.cdl");
import("sTWBasicDispatcherControl.cdl");
import("sTWBasicDispatcherDriverControl.cdl");
import("sTWBasicDispatcherDriverEvent.cdl");
import("sTWDeferredDispatchControl.cdl");
import("tTWDeferredDispatch.cdl");

/** @internal */
[active]
celltype tTWBasicDispatcherCore
{
    entry sTWDispatcherControl eDispatcher;
    entry sTWDispatcherLink eDispatcherLink;
    call sTWTimerManagerLink cTimerManager;
    entry sTWBasicDispatcherControl eBasicDispatcher;
    [optional] call sTWBasicDispatcherDriverControl cDriverControl;
    entry sTWBasicDispatcherDriverEvent eDriverEvent;

    call sTWDeferredDispatchControl cTimeoutDispatch;
    entry sTWDispatchTarget eTimeoutDispatch;

    [optional, dynamic] call sTWDispatchTarget cTarget;

    var {
        intptr_t currentTimeoutToken;
        uint8_t deferredDispatchPending = 0;
    };
};

/**
 * ベアメタル (OS無し) 向けのディスパッチャです。
 */
 [active]
composite tTWBasicDispatcher
{
    /**
     * ディスパッチャの制御に使用する受け口です。
     */
    entry sTWDispatcherControl eDispatcher;

    /**
     * `tTWTimerManager::cDispatcherLink` に結合して下さい。
     */
    entry sTWDispatcherLink eDispatcherLink;

    /**
     * `tTWTimerManager::eTimerManager` に結合して下さい。
     */
    call sTWTimerManagerLink cTimerManager;

    /**
     * `tTWBasicDispatcher` 固有の制御に使用する受け口です。
     */
    entry sTWBasicDispatcherControl eBasicDispatcher;

    /**
     * `tTWBasicDispatcher` のハードウェア依存処理の処理を実装するドライバに結合するための呼び口です。
     */
    [optional] call sTWBasicDispatcherDriverControl cDriverControl;

    /**
     * `tTWBasicDispatcher` のハードウェア依存処理の処理を実装するドライバに結合するための受け口です。
     */
    entry sTWBasicDispatcherDriverEvent eDriverEvent;

    cell tTWDeferredDispatch TimeoutDispatch {
        cTimerManager => composite.cTimerManager;
    };

    cell tTWBasicDispatcherCore Core {
        cTimerManager => composite.cTimerManager;
        cDriverControl => composite.cDriverControl;

        cTimeoutDispatch = TimeoutDispatch.eDeferredDispatch;
        eTimeoutDispatch <= TimeoutDispatch.cTarget;
    };

    eDispatcher => Core.eDispatcher;
    eDispatcherLink => Core.eDispatcherLink;
    eBasicDispatcher => Core.eBasicDispatcher;
    eDriverEvent => Core.eDriverEvent;
};