/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

signature sTWMouseEvent
{
	void mouseDown([in] TWPoint point, [in] uint8_t button);
	void mouseMove([in] TWPoint point);
	void mouseUp([in] TWPoint point, [in] uint8_t button);
};
