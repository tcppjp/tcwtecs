/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTypes.cdl");

/**
 * TCWTecs infrastructure. Do not call any members in the user application.
 * @internal
 */
signature sTWDispatcherLink {
    /**
     * GUIスレッドで、ディスパッチャの `sTWTimerManagerLink::handleDeferredDispatch` を呼出します。
     * `sTWTimerManagerLink::handleDeferredDispatch` の呼出しが行われる前に、これが複数回呼び出されても、
     * `sTWTimerManagerLink::handleDeferredDispatch` がその回数分呼び出される必要はなく、少なくとも1回呼び出される
     * ことのみが保証されます。
     *
     * tTWTimerManager のみがこれを呼出します。
     *
     * `sTWDispatcherControl::invoke` と似ていますが、呼出しは非同期です (`sTWTimerManagerLink::handleDeferredDispatch`
     * の呼出しが完了する前に返ります)。
     *
     * クリティカルセクション内で呼び出されます。
     */
    void startDeferredDispatch(void);

    /**
     * 指定時間後に、ディスパッチャの sTWTimerManagerLink::handleTimeout を呼出します。
     *
     * tTWTimerManager のみがこれを呼出します。
     */
    void setTimeout([in] TWDuration duration);

    /**
     * setTimeout の設定を取り消します。
     *
     * tTWTimerManager のみがこれを呼出します。
     */
    void clearTimeout(void);

    /**
     * クリティカルセクションの開始を要求します。クリティカルセクション中では、アプリケーションは (いかなるコンテクストにおいても)
     * `tTWDeferredDispatch::eDeferredDispatch` への呼出しは行なえません。
     *
     * クリティカルセクションは再帰的であっても良いですが、そうでなくても問題ありません。
     *
     * tTWTimerManager のみがこれを呼出します。
     */
    void enterCriticalSection(void);

    /**
     * クリティカルセクションの終了を要求します。
     *
     * tTWTimerManager のみがこれを呼出します。
     */
    void leaveCriticalSection(void);

    /**
     * 時刻を取得します。基準とする時刻は任意ですが、それは変化してはいけません。また、取得される時刻は stable である必要があります。
     *
     * tTWTimerManager のみがこれを呼出します。
     *
     * @internal
     */
    TWTimePoint getTime(void);
};
