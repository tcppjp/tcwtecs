/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");

signature sTWTimerControl
{
    void setTimeout([in] TWDuration duration, [in] intptr_t param);
    void setInterval([in] TWDuration interval, [in] intptr_t param);
    void clear(void);
};
