/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");
import("sTWDeferredDispatchControl.cdl");
import("sTWTimerManagerLink.cdl");
import("sTWDispatcherControl.cdl");
import("sTWDispatchTarget.cdl");

import_C("TWPrivate.h");

/**
 * Thread-safe mechanism to perform asynchronous dispatch.
 */
celltype tTWDeferredDispatch
{
    entry sTWDeferredDispatchControl eDeferredDispatch;
    call  sTWDispatchTarget          cTarget;

    call sTWTimerManagerLink cTimerManager;

    var {
        TWDeferredDispatchDescriptor descriptor;
    };
};
