/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("tTWView.cdl");
import("tTWDesktop.cdl");
import("tTWTimerManager.cdl");
import("tTWSDLGraphicsDevice.cdl");
import("tTWSDLDispatcher.cdl");
import("tTWKeyboardInputManager.cdl");
import("tTWTouchInputManager.cdl");
import("tTWStaticRectSource.cdl");
import("tTWStaticViewStyleSource.cdl");
