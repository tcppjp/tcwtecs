/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import_C("tecsui/types.h");
import_C("tecsui/geometry.h");
import_C("tecsui/bitmap.h");
import_C("tecsui/colors.h");
