/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("sTWTouchInputDriverEvent.cdl");
import("sTWTouchInputSubviewLink.cdl");
import("sTWTouchInputSuperviewLink.cdl");
import("sTWTouchInputElementLink.cdl");
import_C("tecsui/geometry.h");

/** @private */
celltype tTWTouchInputManagerCore
{
    /** Join this to the root view's `tTWTouchInputElement`'s eSuperview */
    call sTWTouchInputSubviewLink cSubview;

    /** Join this to the root view's `tTWTouchInputElement`'s cSuperview */
    entry sTWTouchInputSuperviewLink eSubview;

    entry sTWTouchInputDriverEvent eDriverEvent;

    attr {
        uint8_t maxNumTouches = 1;
    };

    [dynamic, ref_desc] call sTWTouchInputElementLink cElement[];

    [ref_desc] call sTWTouchInputElementLink cNullElementLink;

    entry sTWTouchInputElementLink eNullElementLink;

    var {
        /**
         * Element-local touch identifiers.
         *
         * WARNING: The value is offseted by one; zero means "nil", and one means
         *          zero (the first touch identifier).
         */
        [size_is(maxNumTouches)] uint8_t *localTouchId;
    };
};

composite tTWTouchInputManager
{
    /** Join this to the root view's `tTWTouchInputElement` */
    call sTWTouchInputSubviewLink cSubview;

    /** Join this to the root view's `tTWTouchInputElement`'s cSuperview */
    entry sTWTouchInputSuperviewLink eSubview;

    entry sTWTouchInputDriverEvent eDriverEvent;

    attr {
        uint8_t maxNumTouches = 1;
    };

    /**
     * This call port array has the number of elements that must much the value
     * of the attribute `maxNumTouches`, and every element should be joined to
     * `eNullElementLink` of the same cell.
     */
    [dynamic, ref_desc] call sTWTouchInputElementLink cElement[];
    entry sTWTouchInputElementLink eNullElementLink;

    cell tTWTouchInputManagerCore Core
    {
        cSubview => composite.cSubview;
        cElement => composite.cElement;
        maxNumTouches = composite.maxNumTouches;

        cNullElementLink = Core.eNullElementLink;
    };

    composite.eSubview => Core.eSubview;
    composite.eDriverEvent => Core.eDriverEvent;
    composite.eNullElementLink => Core.eNullElementLink;
};
