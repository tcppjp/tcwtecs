/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

celltype tTWTouchInputManager
{
    // TODO: tTWTouchInputManager
};
