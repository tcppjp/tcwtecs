/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("sTWTimerManagerLink.cdl");
import("sTWDispatcherLink.cdl");

import_C("TWPrivate.h");

celltype tTWTimerManager
{
    entry sTWTimerManagerLink eTimerManager;

    call sTWDispatcherLink cDispatcherLink;

    var {
        TWPQHeader timerQueue;
        TWDLLHeader timerPendingList;
        TWDLLHeader deferredDispatchQueue;
        uint8_t isProcessingTimers;
    };
};
