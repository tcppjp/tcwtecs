/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import_C("TWSDL2.h");

/**
 * SDLイベントシステムにおけるイベントの伝達に用いられるシグニチャ。
 */
[deviate, callback]
signature sTWSDLEvent
{
    /**
     * SDLイベントシステムのイベントキューにあるイベントを処理する。
     *
     * @return 処理できた場合は 0 以外を返す。処理できなかった場合は 0 を返す。
     */
    uint8_t handle([inout] SDL_Event *event);
};
