/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

/*
 *  This CDL application is well-organized using composite celltypes, but
 *  doesn't work yet with the latest version (at the time of writing) of tecsgen.
 */

import("TWTecs.cdl");

import("tSimpleButton.cdl");

cell tTWSDLGraphicsDevice SDL {
	width = 120;
	height = 120;
	title = "Hello World!";
	windowFlags = C_EXP("0");
};

cell tTWDesktop Desktop {
	cGraphicsDevice = SDL.eGraphicsDevice;
	eGraphicsDevice <= SDL.cGraphicsDevice;
};

celltype tMainWindowCore {
	entry sTWPaintEvent ePaintEvent;
	call sTWDrawingContext cDC;

	entry sAction eButtonActivated[3];
};

composite tMainWindow {
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;
	call sTWDesktopLink cDesktopLink;

	cell tSimpleButton Button1;
	cell tSimpleButton Button2;
	cell tSimpleButton Button3;

	cell tMainWindowCore Core;

	cell tTWStaticRectSource View_Bounds {
		x = 0; y = 0; w = 120; h = 120;
	};
	cell tTWStaticViewStyleSource View_Style {
		value = C_EXP("TWViewStyleVisible");
	};

	cell tTWView View {
		cSuperview => composite.cSuperview;
		cDesktopLink => composite.cDesktopLink;

		cBoundsSource = View_Bounds.eSource;
		cStyleSource = View_Style.eSource;

		// TODO: コールバック結合で記述したい
		cSubview[0] = Button1.eSuperview;
		cSubview[1] = Button2.eSuperview;
		cSubview[2] = Button3.eSuperview;

		cPaintEvent = Core.ePaintEvent;
	};
	composite.eSuperview => View.eSuperview;

	cell tMainWindowCore Core {
		cDC = View.eDrawingContext;
	};

	cell tTWStaticRectSource Button1_Bounds {
		x = 20; y = 20; w = 80; h = 20;
	};
	cell tTWStaticRectSource Button2_Bounds {
		x = 20; y = 50; w = 80; h = 20;
	};
	cell tTWStaticRectSource Button3_Bounds {
		x = 20; y = 80; w = 80; h = 20;
	};
	cell tTWStaticViewStyleSource Button_Style {
		value = C_EXP("TWViewStyleVisible");
	};
	cell tSimpleButton Button1 {
		cSuperview = View.eSubview[0];

		cDesktopLink => composite.cDesktopLink;

		cBoundsSource = Button1_Bounds.eSource;
		cStyleSource = Button_Style.eSource;
		
		cAction = Core.eButtonActivated[0];
	};
	/* TODO: @@cloned_cell_list が同じ複合セルタイプ由来の複数のセルを区別できない問題
	      があるため，tSimpleButton を複数個定義してしまうと結合先がおかしくなる． */
	cell tSimpleButton Button2 {
		cSuperview = View.eSubview[1];

		cDesktopLink => composite.cDesktopLink;

		cBoundsSource = Button2_Bounds.eSource;
		cStyleSource = Button_Style.eSource;
		
		cAction = Core.eButtonActivated[1];
	};
	cell tSimpleButton Button3 {
		cSuperview = View.eSubview[2];

		cDesktopLink => composite.cDesktopLink;

		cBoundsSource = Button3_Bounds.eSource;
		cStyleSource = Button_Style.eSource;
		
		cAction = Core.eButtonActivated[2];
	};
};

cell tMainWindow MainWindow {
	cSuperview = Desktop.eSubview;
	eSuperview <= Desktop.cSubview;
	cDesktopLink = Desktop.eDesktopLink;
};

[active, singleton]
celltype tTestApp {
	call sTWSDLGraphicsDeviceControl cSDL;
	entry sTWSDLGraphicsDeviceEvent eSDL;

	call sTWDesktopControl cDesktop;
};

cell tTestApp App {
	cSDL = SDL.eControl;
	eSDL <= SDL.cEvent;

	cDesktop = Desktop.eDesktop;
};
