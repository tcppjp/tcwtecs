/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTecs.cdl");
import("sAction.cdl");

celltype tSimpleButtonCore {
	entry sTWPaintEvent ePaintEvent;
	entry sTWTouchEvent eTouchEvent;

	// TODO: 本当は optional でいいけど、そうすると composite の非 optional な
	//       call に接続できなくなってしまう! (tecsgen v1.4.0)
	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	call sTWRectSource cBoundsSource;
	call sTWDrawingContext cDrawingContext;
	call sTWViewControl cViewControl;

	[optional] call sAction cAction;

	entry sTWKeyboardEvent eKeyboardEvent;
	[ref_desc] call sTWKeyboardEvent cKeyboardEvent;

	var {
		uint8_t active = 0;
	};
};

composite tSimpleButton {
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;
	call sTWDesktopLink cDesktopLink;

	entry sTWTouchInputSubviewLink eTouchInputSuperview;
	call sTWTouchInputSuperviewLink cTouchInputSuperview;

	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	call sTWViewStyleSource cStyleSource;
	entry sTWValueSourceCallback eStyleSource;

	call sTWRectSource cBoundsSource;
	entry sTWValueSourceCallback eBoundsSource;

	[optional] call sAction cAction;

	cell tSimpleButtonCore Core;
	cell tTWView View;

	cell tSimpleButtonCore Core {
		cBoundsSource => composite.cBoundsSource;
		cAction => composite.cAction;
		cKeyboardInputManager => composite.cKeyboardInputManager;
		cDrawingContext = View.eDrawingContext;
		cViewControl = View.eControl;
		cKeyboardEvent = Core.eKeyboardEvent;
	};

	cell tTWView View {
		cSuperview => composite.cSuperview;
		cDesktopLink => composite.cDesktopLink;

		cBoundsSource => composite.cBoundsSource;
		cStyleSource => composite.cStyleSource;

		cPaintEvent = Core.ePaintEvent;
	};

	cell tTWTouchInputElement TouchInputElement {
		cSuperview => composite.cTouchInputSuperview;

		cTouchEvent = Core.eTouchEvent;

		cBoundsSource => composite.cBoundsSource;
		cStyleSource => composite.cStyleSource;
	};

	cell tTWValueSourceCallbackSplitter BoundsSplitter {
		cCallback[0] = View.eBoundsSource;
		cCallback[1] = TouchInputElement.eBoundsSource;
	};

	cell tTWValueSourceCallbackSplitter StyleSplitter {
		cCallback[0] = View.eStyleSource;
		cCallback[1] = TouchInputElement.eStyleSource;
	};

	composite.eSuperview => View.eSuperview;
	composite.eStyleSource => BoundsSplitter.eCallback;
	composite.eBoundsSource => StyleSplitter.eCallback;
	composite.eTouchInputSuperview => TouchInputElement.eSuperview;
};
