/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");

signature sTWViewControl
{
	TWViewStyle getStyle(void);

	void getBounds([out] TWRect *outRect);
	void getGlobalBounds([out] TWRect *outRect);

	void setNeedsUpdate(void);

	void setFocus(void);
	bool isFocused(void);

	void setMouseCapture(void);
	void releaseMouseCapture(void);
	bool hasMouseCapture(void);
};
