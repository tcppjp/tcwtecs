/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("sTWKeyboardEvent.cdl");

signature sTWKeyboardInputDriverEvent
{
    void notifyKeyDown([in] uint16_t keyCode);
    void notifyKeyUp([in] uint16_t keyCode);
};
