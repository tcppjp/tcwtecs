/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTypes.cdl");
import("sTWSubviewLink.cdl");
import("sTWSuperviewLink.cdl");
import("sTWDesktopLink.cdl");
import("sTWGraphicsDeviceInput.cdl");
import("sTWGraphicsDeviceOutput.cdl");
import("sTWDesktopControl.cdl");

celltype tTWDesktop
{
	entry sTWDesktopControl eDesktop;

	// Join these to the root view
	[optional] call sTWSubviewLink cSubview;
	entry sTWSuperviewLink eSubview;

	// Join these to all views
	entry sTWDesktopLink eDesktopLink;

	// Join to the graphics device
	entry sTWGraphicsDeviceInput eGraphicsDevice;
	call sTWGraphicsDeviceOutput cGraphicsDevice;

	var {
		TWRect dirtyRect;
		TWPoint paintOffset;
	};
};
