/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTecs.cdl");
import("sBitmapData.cdl");

celltype tBitmapViewCore {
    entry sTWPaintEvent ePaintEvent;

    call sTWRectSource cBoundsSource;
    call sTWDrawingContext cDrawingContext;
    call sTWViewControl cViewControl;

    call sBitmapData cBitmapData;
};

composite tBitmapView {
    [optional] call sTWSuperviewLink cSuperview;
    entry sTWSubviewLink eSuperview;
    call sTWDesktopLink cDesktopLink;

    call sTWViewStyleSource cStyleSource;
    entry sTWValueSourceCallback eStyleSource;

    call sTWRectSource cBoundsSource;
    entry sTWValueSourceCallback eBoundsSource;

    call sBitmapData cBitmapData;

    cell tBitmapViewCore Core;
    cell tTWView View;

    cell tBitmapViewCore Core {
        cBoundsSource => composite.cBoundsSource;
        cDrawingContext = View.eDrawingContext;
        cViewControl = View.eControl;

        cBitmapData => composite.cBitmapData;
    };

    cell tTWView View {
        cSuperview => composite.cSuperview;
        cDesktopLink => composite.cDesktopLink;

        cBoundsSource => composite.cBoundsSource;
        cStyleSource => composite.cStyleSource;

        cPaintEvent = Core.ePaintEvent;
    };

    composite.eSuperview => View.eSuperview;
    composite.eStyleSource => View.eStyleSource;
    composite.eBoundsSource => View.eBoundsSource;
};
