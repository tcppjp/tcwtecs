/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

// TODO: keyboard event propagation (through the view hierarchy)
signature sTWKeyboardEvent
{
    /**
     * キー押下時に呼び出されます。
     *
     * @param keyCode TODO
     */
	void keyDown([in] uint16_t keyCode);

    /**
     * キー解放時に呼び出されます。
     *
     * @param keyCode TODO
     */
	void keyUp([in] uint16_t keyCode);

    /**
     * キーボードフォーカス取得直後に呼び出されます。
     *
     * 注意: 本呼び出し中にキーボードフォーカス対象を変更する操作は現時点では未定義動作となります。
     */
    void enter(void);

    /**
     * キーボードフォーカス喪失直前に呼び出されます。
     *
     * 注意: 本呼び出し中にキーボードフォーカス対象を変更する操作は現時点では未定義動作となります。
     */
    void leave(void);
};
