/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("sTWDispatcherControl.cdl");
import("sTWDispatcherLink.cdl");
import("sTWDispatchTarget.cdl");
import("sTWTimerManagerLink.cdl");
import("TWTecs.cdl");

/** @internal */
[singleton, active]
celltype tMyDispatcherCore
{
    entry sTWDispatcherControl eDispatcher;
    entry sTWDispatcherLink eDispatcherLink;
    call sTWTimerManagerLink cTimerManager;
    [optional] call sTWDispatchTarget cInitializer[];
    [optional, dynamic] call sTWDispatchTarget cTarget;

    call sTWDeferredDispatchControl cTimerDispatch;
    entry sTWDispatchTarget eTimerDispatch;
};

[singleton, active]
composite tMyDispatcher
{
    /**
     * ディスパッチャとしての機能を提供する受け口。
     */
    entry sTWDispatcherControl eDispatcher;

    /**
     * `tTWTimerManager::cDispatcherLink` と結合して下さい。
     */
    entry sTWDispatcherLink eDispatcherLink;

    /**
     * `tTWTimerManager::eTimerManager` と結合して下さい。
     */
    call sTWTimerManagerLink cTimerManager;

    /**
     * メインループ開始前に呼ばれるディスパッチターゲット
     */
    [optional] call sTWDispatchTarget cInitializer[];

    cell tTWDeferredDispatch TimerDispatch {
        cTimerManager => composite.cTimerManager;
    };

    cell tMyDispatcherCore Core {
        cTimerManager => composite.cTimerManager;
        cInitializer => composite.cInitializer;

        cTimerDispatch = TimerDispatch.eDeferredDispatch;
        eTimerDispatch <= TimerDispatch.cTarget;
    };

    eDispatcher => Core.eDispatcher;
    eDispatcherLink => Core.eDispatcherLink;
};