/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTypes.cdl");
import("sTWSubviewLink.cdl");
import("sTWSuperviewLink.cdl");
import("sTWViewControl.cdl");
import("sTWDesktopLink.cdl");
import("sTWPaintEvent.cdl");
import("sTWViewStyleSource.cdl");
import("sTWRectSource.cdl");
import("sTWValueSourceCallback.cdl");
import("sTWDrawingContext.cdl");

/**
 * ビューは TCW for TECS における GUI の最小管理単位であり、以下の機能を提供します。
 *
 *  - ビュー階層の表現
 *  - 画面上の占有領域 (境界長方形) の定義
 *  - ビューのコンテンツの描画
 *
 * 基本的な使用方法
 * -------------
 *
 * ビューを使用する為には、以下の使用法に従う必要があります。
 *
 * ### 階層の表現
 *
 * `cSuperView`, `eSuperview`, `cSubview`, `eSubview` を使用して、ビューの階層を表現します。
 * `cSuperView`, `eSuperview` をそれぞれ親ビューの `eSubview`, `cSubview` に結合して下さい。
 * また、 `cDesktopLink` をビューが属するデスクトップの `tTWDesktop::eDesktopLink` に結合する必要があります。
 *
 * ### 境界長方形
 *
 * ビューの境界長方形は、`TWRect` を使用して、親ビュー内のビュー座標系で定義されます。
 * `BoundsSource` プロパティ (`cBoundsSource`, `eBoundsSource` のペア) を使用して境界長方形を定義します。
 *
 * ### 再描画イベントの処理
 *
 * `cPaintEvent::paint` が、ビューの再描画が必要になったときに呼ばれるので、独自に定義したセルにこれを結合してください。
 * これが呼ばれた際には、対応するビューの `eDrawingContext` を経由してビュー全体の描画を行って下さい。
 *
 * `eDrawingContext` の座標系はビューの境界長方形の左上を基準としています。
 *
 * ### ビューの制御
 *
 * `eControl` を呼ぶことにより、ビューの制御が
 *
 * コンポーネント化
 * -------------
 *
 * 新たなタイプのビューを定義する場合、以下のセルを持つ複合セルタイプを定義する必要があります。
 *
 * TODO:
 *
 */
celltype tTWView
{
	// Join these to the superview
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;

	// Join these to subviews
	[optional] call sTWSubviewLink cSubview[];
	entry sTWSuperviewLink eSubview[];

	// Join this to the desktop
	call sTWDesktopLink cDesktopLink;

	// control
	entry sTWViewControl eControl;
	entry sTWDrawingContext eDrawingContext;

	// events
	[optional] call sTWPaintEvent cPaintEvent;

	// properties
	call sTWViewStyleSource cStyleSource;
	entry sTWValueSourceCallback eStyleSource;

	call sTWRectSource cBoundsSource;
	entry sTWValueSourceCallback eBoundsSource;
};
