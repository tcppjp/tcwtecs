/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTecs.cdl");
import("sAction.cdl");

celltype tSimpleButtonCore {
	entry sTWPaintEvent ePaintEvent;
	entry sTWTouchEvent eTouchEvent;

	// TODO: 本当は optional でいいけど、そうすると composite の非 optional な
	//       call に接続できなくなってしまう! (tecsgen v1.4.0)
	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	call sTWRectSource cBoundsSource;
	call sTWDrawingContext cDrawingContext;
	call sTWViewControl cViewControl;

	[optional] call sAction cAction;

	entry sTWKeyboardEvent eKeyboardEvent;
	[ref_desc] call sTWKeyboardEvent cKeyboardEvent;

	var {
		uint8_t active = 0;
	};
};

composite tSimpleButton {
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;
	call sTWDesktopLink cDesktopLink;

	entry sTWTouchInputSubviewLink eTouchInputSuperview;
	call sTWTouchInputSuperviewLink cTouchInputSuperview;

	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	call sTWViewStyleSource cStyleSource;
	entry sTWValueSourceCallback eStyleSource;

	call sTWRectSource cBoundsSource;
	entry sTWValueSourceCallback eBoundsSource;

	[optional] call sAction cAction;

	cell tSimpleButtonCore Core;
	cell tTWView View;

	cell tSimpleButtonCore Core {
		cBoundsSource => composite.cBoundsSource;
		cAction => composite.cAction;
		cKeyboardInputManager => composite.cKeyboardInputManager;
		cDrawingContext = View.eDrawingContext;
		cViewControl = View.eControl;
		cKeyboardEvent = Core.eKeyboardEvent;
	};

	cell tTWView View {
		cSuperview => composite.cSuperview;
		cDesktopLink => composite.cDesktopLink;

		cBoundsSource => composite.cBoundsSource;
		cStyleSource => composite.cStyleSource;

		cPaintEvent = Core.ePaintEvent;
	};

	cell tTWTouchInputElement TouchInputElement {
		cSuperview => composite.cTouchInputSuperview;

		cTouchEvent = Core.eTouchEvent;

		cBoundsSource => composite.cBoundsSource;
		cStyleSource => composite.cStyleSource;
	};

	cell tTWValueSourceCallbackSplitter BoundsSplitter {
		cCallback[0] = View.eBoundsSource;
		cCallback[1] = TouchInputElement.eBoundsSource;
	};

	cell tTWValueSourceCallbackSplitter StyleSplitter {
		cCallback[0] = View.eStyleSource;
		cCallback[1] = TouchInputElement.eStyleSource;
	};

	composite.eSuperview => View.eSuperview;
	composite.eStyleSource => BoundsSplitter.eCallback;
	composite.eBoundsSource => StyleSplitter.eCallback;
	composite.eTouchInputSuperview => TouchInputElement.eSuperview;
};
