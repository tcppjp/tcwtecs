/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");
import("sTWSubviewLink.cdl");
import("sTWSuperviewLink.cdl");
import("sTWDesktopLink.cdl");
import("sTWGraphicsDeviceInput.cdl");
import("sTWGraphicsDeviceOutput.cdl");
import("sTWDesktopControl.cdl");

celltype tTWDesktop
{
	entry sTWDesktopControl eDesktop;

	// Join these to the root view
	[optional] call sTWSubviewLink cSubview;
	entry sTWSuperviewLink eSubview;

	// Join these to all views
	entry sTWDesktopLink eDesktopLink;

	// Join to the graphics device
	entry sTWGraphicsDeviceInput eGraphicsDevice;
	call sTWGraphicsDeviceOutput cGraphicsDevice;

	var {
		void *mouseCaptureTarget = 0;
		void *keyboardFocusTarget = 0;
		TWRect dirtyRect;
		TWPoint paintOffset;
	};
};
