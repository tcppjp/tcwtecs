/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");

[deviate]
signature sTWRenderTargetBitmapSource
{
	void get([out] void **outData, 
		[out] TWPixelFormat *outPixelFormat,
		[out] uint16_t *width, 
		[out] uint16_t *height);
};
