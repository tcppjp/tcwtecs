/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTypes.cdl");

signature sTWDeferredDispatchControl
{
    /**
     * 遅延ディスパッチをスケジュールします。
     *
     * TODO: should update `param` if it's already active?
     *
     * ディスパッチャがクリティカルセクションに進入した状態でない限り、任意のコンテクストから
     * 呼び出せます。
     *
     * @return 既にスケジュール済みであった場合は 0、それ以外の場合は 1。
     */
    uint8_t start([in] intptr_t param);

    /**
     * 遅延ディスパッチをキャンセルします。
     *
     * ディスパッチャがクリティカルセクションに進入した状態でない限り、任意のコンテクストから
     * 呼び出せます。
     *
     * @return スケジュールされていなかった場合は 0、それ以外の場合は 1。
     */
    uint8_t cancel(void);

    // TODO: join (or wait)?
};
