/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");
import("sTWGraphicsDeviceOutput.cdl");
import("sTWRenderTargetBitmapSource.cdl");

import_C("TWPrivate.h");

celltype tTWRGB565BitmapGraphicsRenderer
{
	entry sTWGraphicsDeviceOutput eGraphicsDeviceOutput;
	call sTWRenderTargetBitmapSource cRenderTargetBitmapSource;

    attr {
        uint16_t numScanlineClipperNodes = 256;
    };

	var {
        TWRect scissor;

        TWScanlineClipperState scanlineClipper;
        TWScanlineClipperLineScanState scanlineClipperLineScanner;

        [size_is(numScanlineClipperNodes)]
        TWScanlineClipperNode *scanlineClipperNodes;
	};
};
