/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

signature sTWSDLDispatcherControl
{
    /**
     * SDL2用ディスパッチャを初期化します。
     *
     * この呼出しを行う前に、`SDL_Init` または `SDL_InitSubSystem` を使用し、少なくとも `SDL_INIT_EVENTS`, `SDL_INIT_TIMER`
     * サブシステムの初期化を行う必要があります。
     *
     * 本関数はメインスレッドでのみ呼び出せます。
     */
    void initialize(void);

    /**
     * メインイベントループを開始します。
     *
     * この関数は、`quit()` が呼び出されるか、`SDL_QUIT` イベントが発生するまで返りません。
     *
     * 本関数はメインスレッドでのみ呼び出せます。
     */
    void enterMainLoop(void);

    /**
     * イベントループを抜けさせます。
     *
     * 本関数は任意のスレッドで呼び出せます。
     */
    void quit(void);
};
