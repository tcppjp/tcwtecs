/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("sTWKeyboardEvent.cdl");

signature sTWKeyboardInputManagerControl
{
    void setEventReceiver([in] Descriptor(sTWKeyboardEvent) receiver);
    void clearEventReceiver(void);

    uint8_t isEventReceiver([in] Descriptor(sTWKeyboardEvent) receiver);
};
