/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("sTWKeyboardInputManagerControl.cdl");
import("sTWKeyboardInputDriverEvent.cdl");
import("sTWKeyboardEvent.cdl");

celltype tTWKeyboardInputManager
{
    entry sTWKeyboardInputManagerControl eControl;
    entry sTWKeyboardInputDriverEvent eDriverEvent;

    /** Used internally; do not make any attempt to join this to anything */
    [dynamic, optional, ref_desc] call sTWKeyboardEvent cReceiver;
};
