/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

/**
 * TCWTecs infrastructure. Do not call any members in the user application.
 */
[deviate]
signature sTWDesktopLink
{
	// proxy of sTWDrawingContext
	void fillRect([in] TWColor color, [in] const TWRect *rect);
	void drawBitmap(
		[in, size_is(numBytes)] const char *data,
        [in] uint32_t numBytes,
        [in] const TWBitmapInfo *info,
        [in] uint16_t infoSize,
		[in] const TWRect *inRect,
		[in] const TWPoint *outLoc);
	void preparePaint([in] const TWRect *globalClipRect, [in] const TWPoint *globalLoc);
	void subtractClippingRect([in] const TWRect *globalClipRect);
};
