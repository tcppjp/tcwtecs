/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTecs.cdl");
import("sAction.cdl");

celltype tSimpleButtonCore {
	entry sTWPaintEvent ePaintEvent;
	entry sTWMouseEvent eMouseEvent;
	entry sTWFocusEvent eFocusEvent;

	// TODO: 本当は optional でいいけど、そうすると composite の非 optional な
	//       call に接続できなくなってしまう! (tecsgen v1.4.0)
	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	call sTWRectSource cBoundsSource;
	call sTWDrawingContext cDrawingContext;
	call sTWViewControl cViewControl;

	[optional] call sAction cAction;

	/** 自身の cKeyboardEvent と結合して下さい。 */
	entry sTWKeyboardEvent eKeyboardEvent;
	/** 自身の eKeyboardEvent と結合して下さい。 */
	[ref_desc] call sTWKeyboardEvent cKeyboardEvent;
};

composite tSimpleButton {
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;
	call sTWDesktopLink cDesktopLink;

	call sTWKeyboardInputManagerControl cKeyboardInputManager;

	call sTWViewStyleSource cStyleSource;
	entry sTWValueSourceCallback eStyleSource;

	call sTWRectSource cBoundsSource;
	entry sTWValueSourceCallback eBoundsSource;

	[optional] call sAction cAction;

	cell tSimpleButtonCore Core;
	cell tTWView View;

	cell tSimpleButtonCore Core {
		cBoundsSource => composite.cBoundsSource;
		cAction => composite.cAction;
		cKeyboardInputManager => composite.cKeyboardInputManager;
		cDrawingContext = View.eDrawingContext;
		cViewControl = View.eControl;
		cKeyboardEvent = Core.eKeyboardEvent;
	};

	cell tTWView View {
		cSuperview => composite.cSuperview;
		cDesktopLink => composite.cDesktopLink;

		cBoundsSource => composite.cBoundsSource;
		cStyleSource => composite.cStyleSource;

		cPaintEvent = Core.ePaintEvent;
		cMouseEvent = Core.eMouseEvent;
		cFocusEvent = Core.eFocusEvent;
	};

	composite.eSuperview => View.eSuperview;
	composite.eStyleSource => View.eStyleSource;
	composite.eBoundsSource => View.eBoundsSource;
};
