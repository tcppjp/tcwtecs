/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("sTWDispatcherControl.cdl");
import("sTWDispatcherLink.cdl");
import("sTWDispatchTarget.cdl");
import("sTWTimerManagerLink.cdl");
import("sTWSDLDispatcherControl.cdl");
import("sTWSDLEvent.cdl");

// It's singleton because SDL2 doesn't support multple event queues
[singleton]
celltype tTWSDLDispatcher
{
    /**
     * ディスパッチャとしての機能を提供する受け口。
     */
    entry sTWDispatcherControl eDispatcher;

    /**
     * `tTWSDLDispatcher` に固有の機能を提供する受け口。
     */
    entry sTWSDLDispatcherControl eSDLDispatcher;

    /**
     * `tTWTimerManager::cDispatcherLink` と結合して下さい。
     */
    entry sTWDispatcherLink eDispatcherLink;

    /**
     * `tTWTimerManager::eTimerManager` と結合して下さい。
     */
    call sTWTimerManagerLink cTimerManager;

    /**
     * SDLイベントシステムを利用してイベントを受け取るための呼び口。
     */
    [optional] call sTWSDLEvent cSDLEvent[];

    /**
     * 内部的に使用されます。結合しないで下さい。
     * @internal
     */
    [optional, dynamic] call sTWDispatchTarget cTarget;
};