/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

import("TWTypes.cdl");
import("sTWGraphicsDeviceOutput.cdl");
import("sTWRenderTargetBitmapSource.cdl");

celltype tTWRGBX32BitmapGraphicsRenderer
{
	entry sTWGraphicsDeviceOutput eGraphicsDeviceOutput;
	call sTWRenderTargetBitmapSource cRenderTargetBitmapSource;

	var {
		TWRect scissor;
	};
};
