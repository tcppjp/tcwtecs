/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("TWTypes.cdl");
import("sTWSubviewLink.cdl");
import("sTWSuperviewLink.cdl");
import("sTWViewControl.cdl");
import("sTWDesktopLink.cdl");
import("sTWMouseEvent.cdl");
import("sTWKeyboardEvent.cdl");
import("sTWPaintEvent.cdl");
import("sTWViewStyleSource.cdl");
import("sTWRectSource.cdl");
import("sTWValueSourceCallback.cdl");
import("sTWDrawingContext.cdl");

celltype tTWView
{
	// Join these to the superview
	[optional] call sTWSuperviewLink cSuperview;
	entry sTWSubviewLink eSuperview;

	// Join these to subviews
	[optional] call sTWSubviewLink cSubview[];
	entry sTWSuperviewLink eSubview[];

	// Join this to the desktop
	call sTWDesktopLink cDesktopLink;

	// control
	entry sTWViewControl eControl;
	entry sTWDrawingContext eDrawingContext;

	// events
	[optional] call sTWMouseEvent cMouseEvent;
	[optional] call sTWPaintEvent cPaintEvent;

	// properties
	call sTWViewStyleSource cStyleSource;
	entry sTWValueSourceCallback eStyleSource;

	call sTWRectSource cBoundsSource;
	entry sTWValueSourceCallback eBoundsSource;
};
