/*
 * Copyright (C) 2016 Tomoaki Kawada
 *
 * This software may be modified and distributed under the terms
 * of the MIT license.  See the LICENSE file for details.
 */

/** 
 * TCWTecs infrastructure. Do not call any members in the user application.
 */
[deviate]
signature sTWDesktopLink
{
	// focus management
	void *getMouseCaptureTarget(void);
	void setMouseCaptureTarget([inout] void *newTarget);

	// proxy of sTWDrawingContext
	void fillRect([in] TWColor color, [in] const TWRect *rect);
	void drawBitmap(
		[in, size_is(numBytes)] const char *data, 
		[in] TWPixelFormat format,
		[in] const TWSize *bitmapSize,
		[in] uint32_t numBytes,
		[in] const TWRect *inRect,
		[in] const TWPoint *outLoc,
		[in] TWColor monoColor);
	void preparePaint([in] const TWRect *globalClipRect, [in] const TWPoint *globalLoc);
};
