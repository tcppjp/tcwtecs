/*
 * Copyright (C) 2017 Tomoaki Kawada
 *
 * This file is part of tcwtecs.
 *
 * tcwtecs is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * tcwtecs is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with tcwtecs.  If not, see <http://www.gnu.org/licenses/>.
 */

import("sTWGraphicsDeviceInput.cdl");
import("sTWGraphicsDeviceOutput.cdl");
import("tTWRGBX32BitmapGraphicsRenderer.cdl");
import("sTWSDLGraphicsDeviceControl.cdl");
import("sTWSDLEvent.cdl");
import("sTWKeyboardInputDriverEvent.cdl");
import("sTWTouchInputDriverEvent.cdl");

/** @internal */
celltype tTWSDLGraphicsDeviceCore
{
	entry sTWRenderTargetBitmapSource eBitmapSource;

	entry sTWGraphicsDeviceOutput eOutput;
	call sTWGraphicsDeviceOutput cOutput;

	call sTWKeyboardInputDriverEvent cKeyboardInputDriverEvent;
	call sTWTouchInputDriverEvent cTouchInputDriverEvent;

	entry sTWSDLGraphicsDeviceControl eControl;

	entry sTWSDLEvent eSDLEvent; // TODO: implement this!

	attr {
		uint16_t width;
		uint16_t height;
		const char *title;
		uint32_t windowFlags;
	};

	var {
		void *window;
		void *surface;
	};
};

/**
 * Example implementation of graphics device for SDL (Simple DirectMedia Library).
 */
composite tTWSDLGraphicsDevice
{
	call sTWKeyboardInputDriverEvent cKeyboardInputDriverEvent;
	call sTWTouchInputDriverEvent cTouchInputDriverEvent;
	entry sTWGraphicsDeviceOutput eGraphicsDevice;

	entry sTWSDLGraphicsDeviceControl eControl;

	entry sTWSDLEvent eSDLEvent;

	attr {
		uint16_t width;
		uint16_t height;
		const char *title;
		uint32_t windowFlags;
	};

	cell tTWSDLGraphicsDeviceCore Core;
	cell tTWRGBX32BitmapGraphicsRenderer Renderer;

	cell tTWSDLGraphicsDeviceCore Core {
		cKeyboardInputDriverEvent => composite.cKeyboardInputDriverEvent;
		cTouchInputDriverEvent => composite.cTouchInputDriverEvent;
		width = composite.width;
		height = composite.height;
		title = composite.title;
		windowFlags = composite.windowFlags;
		cOutput = Renderer.eGraphicsDeviceOutput;
	};
	cell tTWRGBX32BitmapGraphicsRenderer Renderer {
		cRenderTargetBitmapSource = Core.eBitmapSource;
	};

	eGraphicsDevice => Core.eOutput;
	eControl => Core.eControl;
	eSDLEvent => Core.eSDLEvent;
};
